`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.10.2022 17:13:07
// Design Name: 
// Module Name: DDL4x4Luma
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module DDR4x4Luma(
    input clk,
    input reset,
    input [7:0] A,
    input [7:0] B,
    input [7:0] C,
    input [7:0] D,
    input [7:0] E,
    input [7:0] F,
    input [7:0] G,
    input [7:0] H,
    input [7:0] I,
    input [7:0] J,
    input [7:0] K,
    input [7:0] L,
    input [7:0] M,
    output reg [7:0] ddrpred [15:0]
    );
    
        always @(posedge clk) begin
            ddrpred[0] <= (I+2*M+A+2)>>2; //a
            ddrpred[1] <= (M+2*A+B+2)>>2;//b
            ddrpred[2] <= (A+2*B+C+2)>>2;//c
            ddrpred[3] <= (B+2*C+D+2)>>2;//d
            ddrpred[4] <= (J+2*I+M+2)>>2;//e
            ddrpred[5] <= (I+2*M+A+2)>>2;//f
            ddrpred[6] <= (M+2*A+B+2)>>2;//g
            ddrpred[7] <= (A+2*B+C+2)>>2;//h
            ddrpred[8] <= (K+2*J+I+2)>>2;//i
            ddrpred[9] <= (J+2*I+M+2)>>2;//j
            ddrpred[10] <=(I+2*M+A+2)>>2;//k
            ddrpred[11] <=(M+2*A+B+2)>>2;//l
            ddrpred[12] <=(L+2*K+J+2)>>1;//m
            ddrpred[13] <=(K+2*J+I+2)>>2;//n
            ddrpred[14] <=(J+2*I+M+2)>>2;//o
            ddrpred[15] <=(I+2*M+A+2)>>2;//[       
        end     
        

endmodule